MemoriaTeste_inst : MemoriaTeste PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
