library verilog;
use verilog.vl_types.all;
entity processadorSch_vlg_vec_tst is
end processadorSch_vlg_vec_tst;
